`define      Idle     3'b001
`define      Start    3'b010
`define      Data     3'b011
`define      Stop     3'b100

    
`define               Display_zero                7'h30
`define               Display_one                 7'h79   
`define               Display_two                 7'h24  
`define               Display_three               7'h30

`define               Display_four                7'h19    
`define               Display_five                7'h12    
`define               Display_six                 7'h2     
`define               Display_seven               7'h78
 
`define               Display_eight               7'h0 
`define               Display_nine                7'h6f
`define               Display_a                   7'h1f
